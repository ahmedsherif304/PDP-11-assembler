library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

Entity ROM is
port (
clk : in std_logic;
uAR : in std_logic_vector(8 downto 0);
CW : out std_logic_vector(31 downto 0) );
end entity ROM;

architecture ROM_Arc of ROM is
	type ROM_type is array(0 to 512) of std_logic_vector(31 downto 0);

	signal rom : ROM_type := (
0   	=>  	"00000000100101101000101011100000",
1   	=>  	"00000001001100100000000000010000",
2   	=>  	"00000000001001000000000000000001",
3   	=>  	"00000100000000000000000000000000",
4	=>	"00000000000000000000000000000000",
5 	=> 	"00000011000100000010000000000000",
6	=> 	"00000011100001100010100000000001",
7	=> 	"00000000001100100000000000000000",
65	=>	"01000000110000000100000000000010",
73	=>	"00111011110000001000000010000000",
81	=>	"00101001010001101000101011100000",
82	=>	"00111011001110000000000000010100",
97	=>	"00110001010001101000111011100000",
98	=>	"00111011001110000000000000010100",
113	=>	"00111001000101101000101011100000",
114	=>	"00111001101100100000000000000000",
115	=>	"00111010010000000010000000010000",
116	=>	"00111010101001100000100000000000",
117	=>	"00111011001100001000000010010100",
118	=>	"00111011101000001000000010010000",
119	=>	"01000000101000000100000000000010",
129	=>	"01100001110100000110000000001110",
137	=>	"01011011110100001000000010010000",
145	=>	"01001001010101101000101011100000",
146	=>	"01011011001110100000000000010110",
161	=>	"01010001010101101000111011100000",
162	=>	"01011011001110100000000000010110",
177	=>	"01011001000101101000101011100000",
178	=>	"01011001101100100000000000000000",
179	=>	"01011010010100000010000000010000",
180	=>	"01011010101001100000100000000000",
181	=>	"01011011001100001000000010010110",
182	=>	"01011011101000001000000010010000",
183	=>	"01100001101000000110000000001110",
186	=>	"00000000001100010000000100010000",
187	=>	"00000000001100000110000000000000",
195     =>      "01011101011001100000100001001000",
196     =>      "10001000011000000010000000000000",
272     =>      "01011101011101100000100000001000",
197     =>      "10001000111000000010000000000000",
273     =>      "01011101011101100000101000001000",
198     =>      "10001001011000000010000000000000",
274     =>      "01011101011101100000110000001000",
199     =>      "10001001111000000010000000000000",
275     =>      "01011101011101100000111000001000",
200     =>      "10001010011000000010000000000000",
276     =>      "01011101011101100001000000001000",
201     =>      "10001010111000000010000000000000",
277     =>      "01011101011101100001001000001000",
202     =>      "10001011011000000010000000000000",
278     =>      "01011101011101100001010000001000",
203     =>      "10001011111000000010000000000000",
279     =>      "00000000011101100001011000000000",
259     =>      "01011101011101100000101001101000",
260     =>      "01011101011101100000111001101000",
261     =>      "01011101011101100010110000001000",
262     =>      "01011101011101100000001000001000",
263     =>      "01011101011101100000010000001000",
264     =>      "01011101011101100000011000001000",
265     =>      "01011101011101100001100000001000",
266     =>      "01011101011101100001101000001000",
267     =>      "01011101011101100001110000001000",
others => "00000000000000000000000000000000"
);-- if next address is 10 then end the program
	begin
		process(clk) is
		  Begin
			if rising_edge(clk) then  
				CW <= rom(to_integer(unsigned(uAR)));
			end if;
		end process;

end architecture ROM_Arc;