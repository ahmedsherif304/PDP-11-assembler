library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

Entity ROM is
port (
clk : in std_logic;
uAR : in std_logic_vector(8 downto 0);
CW : out std_logic_vector(31 downto 0) );
end entity ROM;

architecture ROM_Arc of ROM is
	type ROM_type is array(0 to 512) of std_logic_vector(31 downto 0);

	signal rom : ROM_type := (
0   	=>  	"00000000100101101000100011100000",
1   	=>  	"00000001001100100000000000010000",
2   	=>  	"00000000001001000000000000000001",
3   	=>  	"00000100000000000000000000000000",
4	=>	"00000000000000000000000000000000",
5 	=> 	"00000011000100000010000000000000",
6	=> 	"00000011100001100010100000000001",
7	=> 	"00000000001100100000000000000000",
101	=>	"01000000110000000100000000000010",
111	=>	"00111011110000001000000010000000",
121	=>	"00101001010001101000101011100000",
122	=>	"00111011001110000000000000010100",
141	=>	"00110001010001101000111011100000",
142	=>	"00111011001110000000000000010100",
161	=>	"00111001000101101000101011100000",
162	=>	"00111001101100100000000000000000",
163	=>	"00111010010000000010000000010000",
164	=>	"00111010101001100000100000000000",
165	=>	"00111011001100001000000010010100",
166	=>	"00111011101000001000000010010000",
167	=>	"01000000101000000100000000000010",
201	=>	"01100001110100000110000000001110",
211	=>	"01011011110100001000000010010000",
221	=>	"01001001010101101000101011100000",
222	=>	"01011011001110100000000000010110",
241	=>	"01010001010101101000111011100000",
242	=>	"01011011001110100000000000010110",
261	=>	"01011001000101101000101011100000",
262	=>	"01011001101100100000000000000000",
263	=>	"01011010010100000010000000010000",
264	=>	"01011010101001100000100000000000",
265	=>	"01011011001100001000000010010110",
266	=>	"01011011101000001000000010010000",
267	=>	"01100001101000000110000000001110",
272	=>	"00000000001100010000000100010000",
273	=>	"00000000001100000110000000000000",
303     =>      "01011101011001100000100001001000",
304     =>      "10001000011000000010000000000000",
420     =>      "01011101011101100000100000001000",
305     =>      "10001000111000000010000000000000",
421     =>      "01011101011101100000101000001000",
306     =>      "10001001011000000010000000000000",
422     =>      "01011101011101100000110000001000",
307     =>      "10001001111000000010000000000000",
423     =>      "01011101011101100000111000001000",
310     =>      "10001010011000000010000000000000",
424     =>      "01011101011101100001000000001000",
311     =>      "10001010111000000010000000000000",
425     =>      "01011101011101100001001000001000",
312     =>      "10001011011000000010000000000000",
426     =>      "01011101011101100001010000001000",
313     =>      "10001011111000000010000000000000",
427     =>      "00000000011101100001011000000000",
403     =>      "01011101011101100000101001101000",
404     =>      "01011101011101100000111001101000",
405     =>      "01011101011101100010110000001000",
406     =>      "01011101011101100000001000001000",
407     =>      "01011101011101100000010000001000",
410     =>      "01011101011101100000011000001000",
411     =>      "01011101011101100001100000001000",
412     =>      "01011101011101100001101000001000",
413     =>      "01011101011101100001110000001000",
others => "00000000000000000000000000000000"
);-- if next address is 10 then end the program
	begin
		process(clk) is
		  Begin
			if falling_edge(clk) then  
				CW <= rom(to_integer(unsigned(uAR)));
			end if;
		end process;

end architecture ROM_Arc;